//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module arithmetic_right_shift_of_N_by_S_using_arithmetic_right_shift_operation
# (parameter N = 8, S = 3)
(input  [N - 1:0] a, output [N - 1:0] res);

  wire signed [N - 1:0] as = a;
  assign res = as >>> S;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module arithmetic_right_shift_of_N_by_S_using_concatenation
# (parameter N = 8, S = 3)
(input  [N - 1:0] a, output [N - 1:0] res);

  // Task:
  //
  // Implement a module with the logic for the arithmetic right shift,
  // but without using ">>>" operation. You are allowed to use only
  // concatenations ({a, b}), bit repetitions ({ a { b }}), bit slices
  // and constant expressions.

  logic [N - 1:0] shifted_part;
  logic sign_bit;

  assign shifted_part = a[N - 1:0] >> S;
  assign sign_bit = a[N - 1];
  assign res = (S == 0) ? a : (S >= N) ? { N{sign_bit} } : 
                                         { { S{sign_bit} }, shifted_part[N - S - 1:0] };

endmodule

module arithmetic_right_shift_of_N_by_S_using_for_inside_always
# (parameter N = 8, S = 3)
(input  [N - 1:0] a, output logic [N - 1:0] res);

  // Task:
  //
  // Implement a module with the logic for the arithmetic right shift,
  // but without using ">>>" operation, concatenations or bit slices.
  // You are allowed to use only "always_comb" with a "for" loop
  // that iterates through the individual bits of the input.

  always_comb begin
    if (S == 0) begin
      res = a;
    end else if (S >= N) begin
      for (int i = 0; i < N; i++) begin
        res[i] = a[N - 1];
      end
    end else begin
      for (int i = 0; i < N; i++) begin
        if (i + S < N) begin
          res[i] = a[i + S];
        end else begin
          res[i] = a[N - 1];
        end
      end
    end
  end

endmodule

module arithmetic_right_shift_of_N_by_S_using_for_inside_generate
# (parameter N = 8, S = 3)
(input  [N - 1:0] a, output [N - 1:0] res);

  // Task:
  // Implement a module that arithmetically shifts input exactly
  // by `S` bits to the right using "generate" and "for"

  genvar i;
  generate
    for (i = 0; i < N; i = i + 1) begin
      if (i + S < N) begin
        assign res[i] = a[i + S];
      end else begin
        assign res[i] = a[N - 1];
      end
    end
  endgenerate

endmodule
